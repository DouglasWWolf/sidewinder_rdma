
//================================================================================================
//    Date         Version     Who  Changes
// -----------------------------------------------------------------------------------------------
// 25-Oct-2023     1.0.0       DWW  Initial creation
//================================================================================================
localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;

localparam VERSION_DAY   = 25;
localparam VERSION_MONTH = 10;
localparam VERSION_YEAR  = 2023;
